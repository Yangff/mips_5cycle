module alu_decoder(funt, alu_op);
    
endmodule